
`timescale       1ns/1ps


module           testfifo3_3();
    reg                 clk         ; 
    reg                 rst_n       ;
    reg                 din_vld     ;
    reg                 din_sop     ;
    reg       [15:0]    din         ;
    reg                 din_eop     ;
    reg                 din_err     ;       //  Error Package indicator; 
 
    wire                dout_vld    ;
    wire                dout_sop    ;
    wire      [15:0]    dout        ;
    wire                dout_eop    ;  



    parameter   PERIOD    = 20;   // ʱ�����ڣ���λΪns;
    parameter   RST_TIME  = 3 ;   // ��λʱ�䣬��ʱ��ʾ��λ3��ʱ�����ڵ�ʱ�䡣


    integer     i;
    integer     j;


    // ������ģ�������
    fifo_p uut_FIFO_exac_1633(
                                .clk        (   clk        ),        
                                .rst_n      (   rst_n      ),
                                .din_vld    (   din_vld    ),
                                .din_sop    (   din_sop    ),
                                .din        (   din        ),
                                .din_eop    (   din_eop    ),
                                .din_err    (   din_err    ),
                                                         
                                .dout_vld   (   dout_vld   ),
                                .dout_sop   (   dout_sop   ),
                                .dout       (   dout       ),
                                .dout_eop   (   dout_eop   )   
                                );



    //���ɱ���ʱ��50M��Ҳ���� always ���(ͬ��Ҫ�ȶ� clk �� initial ��ʼ����ֵ)��  always  #10  clk = ~clk;
    initial  begin
        clk = 1;
        forever   #(PERIOD/2)    clk=~clk;
    end



    // ������λ�ź�
    initial  begin
        rst_n = 1;
        #2;
        rst_n = 0;
        repeat(3)@(negedge clk);   // ���������� rst_n ��λ�ź�ʱ����ý� clk �ĳ�ʼ��ֵ��Ϊ clk==1��
        rst_n = 1;
    end




    // �����ź�din1��ֵ��ʽ
    initial  begin
        #1;              // ����ֵ
        din_vld = 0;
        din_sop = 0;
        din     = 16'h0;  
        din_eop = 0;
        din_err = 0;     

        #(10*PERIOD);    // ��ʼ��ֵ

        for(j=1; j<4; j=j+1) begin

            for(i=1; i<66; i=i+1) begin
                din_vld =  1;
                din_sop = (i==1)?1:0;
                din     =  i; 
                din_eop = (i==65)?1:0;
                din_err = (i==65 && j==2)?1:0; 
                #(1*PERIOD);
            end 

            din_vld = 0;
            din_sop = 0;
            din     = 16'h0;  
            din_eop = 0;
            din_err = 0;     
            #(10*PERIOD); 
        end
        
        din_vld = 0;
        din_sop = 0;
        din     = 16'h0;  
        din_eop = 0;
        din_err = 0;  

    end




endmodule




